`define OP_LSL 4'h0
`define OP_LSR 4'h1
`define OP_CSL 4'h2
`define OP_CSR 4'h3
`define OP_ASR 4'h4
`define OP_AND 4'h5
`define OP_OR 4'h6
`define OP_XOR 4'h7
`define OP_ADD 4'h8
`define OP_NOP 4'h9
